`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:04:00 11/21/2013 
// Design Name: 
// Module Name:    invsubbyteShiftRow 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module invsubbyteShiftRow(
    input [127:0] in,
    output [127:0] out
    );
wire [127:0] temp;

invsubbyte s0(.out(temp[127:120]),.in(in[127:120]));        
invsubbyte s1(.out(temp[119:112]),.in(in[119:112]));
invsubbyte s2(.out(temp[111:104]),.in(in[111:104]));
invsubbyte s3(.out(temp[103:96]),.in(in[103:96]));

invsubbyte s4(.out(temp[95:88]),.in(in[95:88]));
invsubbyte s5(.out(temp[87:80]),.in(in[87:80]));
invsubbyte s6(.out(temp[79:72]),.in(in[79:72]));
invsubbyte s7(.out(temp[71:64]),.in(in[71:64]));

invsubbyte s8(.out(temp[63:56]),.in(in[63:56]));
invsubbyte s9(.out(temp[55:48]),.in(in[55:48]));
invsubbyte s10(.out(temp[47:40]),.in(in[47:40]));
invsubbyte s11(.out(temp[39:32]),.in(in[39:32]));

invsubbyte s12(.out(temp[31:24]),.in(in[31:24]));
invsubbyte s13(.out(temp[23:16]),.in(in[23:16]));
invsubbyte s14(.out(temp[15:8]),.in(in[15:8]));
invsubbyte s15(.out(temp[7:0]),.in(in[7:0]));

invshiftRow R1(.in(temp),.out(out));

endmodule
